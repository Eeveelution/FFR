module control (
    input wire clk
);


endmodule